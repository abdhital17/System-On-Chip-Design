module brd(
    input clk,
    input enable,
    input [23:0] ibrd,
    input [7:0] fbrd,
    output out
    );
    
endmodule